module data_mem(
	input clk,
	input []addr,
	input []data_in,
	input []op,
	input we,
	output data_out
);

endmodule
