module instr_mem(
	input []addr;
	output []data
);

endmodule
