module cpu(
	input clk,
	input rst
);

endmodule
